module IFU #(DATA_WIDTH = 32) (
  input clk,
  input rst,
  input [DATA_WIDTH-1:0] pc
  //output reg [DATA_WIDTH-1:0] pc_d,
);

  always @(posedge clk) begin
    if (!rst) begin

    end
    else begin 

    end
  end
  
endmodule
