module IFU #(DATA_WIDTH = 32) (
  input clk,
  input rst,
  input [DATA_WIDTH-1:0] pc,
  output reg [DATA_WIDTH-1:0] inst
);

  
endmodule
